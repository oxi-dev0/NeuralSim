CIRCLE 0 64 25
CIRCLE 128 64 25