IF {STEP} > 75
BOX 64 128 0 128
ELSE
CIRCLE 64 64 25
ENDIF